library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity schaltung_b is
  port ( A : in  std_logic;
         B : in  std_logic;
         C : in  std_logic;
         D : in  std_logic;
         Y : out std_logic);
end schaltung_b;

architecture Behavioral of schaltung_b is

begin
  --Direkte zuweisung der Funktion auf
  --den Ausgang

end Behavioral;


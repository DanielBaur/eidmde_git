library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity KV_b is
  port ( --Ein und Ausgaenge definieren
  );
end KV_b;

architecture Behavioral of KV_b is

begin
 --OUT<= minimaler disjunktiver Ausdruck;
end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity KV_a is
  port (
  --Ein und Ausgaenge definieren
  );
end KV_a;

architecture Behavioral of KV_a is

begin

--OUT<= Disjunktive Normalform;
		
end Behavioral;


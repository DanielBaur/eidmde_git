
-- ----------------------------------------
-- libraries
-- ----------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



-- ----------------------------------------
-- entity
-- ----------------------------------------

entity and_gate is
    Port (

        -- Define input and output signals here.

    );
end and_gate;



-- ----------------------------------------
-- architecture
-- ----------------------------------------

architecture Behavioral of and_gate is

begin

    -- Assign signals here.

end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity and_gate is
    Port ( 
           --hier Signale definieren in:A,B; out C
           );
end and_gate;

architecture Behavioral of and_gate is

begin
--Zuweisung C<=?


end Behavioral;


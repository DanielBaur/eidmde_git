library IEEE;
use IEEE.STD_LOGIC_1164.all;

Library UNISIM;
use UNISIM.vcomponents.all;

entity KV_c is
  port ( --Ein und Ausgaenge definieren
  );
end KV_c;

architecture Behavioral of KV_c is



begin

--LUT4_L instanzieren (siehe edit/Language Templates/VHDL/Device Primitive Instatiation/Spartan3/Slice CLB Primitives/LUTs/LUT4_L)
--und init setzen (siehe edit/Language Templates/VHDL/Device Primitive Instatiation/Spartan3/Slice CLB Primitives/LUTs/Info)
--+ Verbindungen mit Ein und Ausgaengen 



end Behavioral;
